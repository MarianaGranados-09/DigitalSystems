library IEEE;
use IEEE.STD_LOGIC_1164.ALL;  

Entity SineLUT is 
	port(
	ANG: in std_logic_vector(6 downto 0);
	SIN: out std_logic_vector(10 downto 0)
);
end SineLUT;

Architecture DataFlow of SineLUT is
begin
	With ANG select SIN <=
	  	--"00000000000" when "0000000",
		"00010010011" when "0000001",
		"00100100110" when "0000010",
		"00110111000" when "0000011",
		"01001001001" when "0000100",
		"01011011000" when "0000101",
		"01101100110" when "0000110",
		"01111110010" when "0000111",
		"10001111100" when "0001000",
		"10100000010" when "0001001",
		"10110000110" when "0001010",
		"11000000110" when "0001011",
		"11010000010" when "0001100",
		"11011111011" when "0001101",
		"11101101111" when "0001110",
		"11111011110" when "0001111",
		"00001001001" when "0010000",
		"00010101110" when "0010001",
		"00100001111" when "0010010",
		"00101101001" when "0010011",
		"00110111110" when "0010100",
		"01000001101" when "0010101",
		"01001010101" when "0010110",
		"01010010111" when "0010111",
		"01011010011" when "0011000",
		"01100001000" when "0011001",
		"01100110110" when "0011010",
		"01101011110" when "0011011",
		"01101111110" when "0011100",
		"01110010111" when "0011101",
		"01110101001" when "0011110",
		"01110110100" when "0011111",
		"01110111000" when "0100000",
		"01110110100" when "0100001",
		"01110101001" when "0100010",
		"01110010111" when "0100011",
		"01101111110" when "0100100",
		"01101011110" when "0100101",
		"01100110110" when "0100110",
		"01100001000" when "0100111",
		"01011010011" when "0101000",
		"01010010111" when "0101001",
		"01001010101" when "0101010",
		"01000001101" when "0101011",
		"00110111110" when "0101100",
		"00101101001" when "0101101",
		"00100001111" when "0101110",
		"00010101110" when "0101111",
		"00001001001" when "0110000",
		"11111011110" when "0110001",
		"11101101111" when "0110010",
		"11011111011" when "0110011",
		"11010000010" when "0110100",
		"11000000110" when "0110101",
		"10110000110" when "0110110",
		"10100000010" when "0110111",
		"10001111100" when "0111000",
		"01111110010" when "0111001",
		"01101100110" when "0111010",
		"01011011000" when "0111011",
		"01001001001" when "0111100",
		"00110111000" when "0111101",
		"00100100110" when "0111110",
		"00010010011" when "0111111",
		"00000000000" when "1000000",
		"00010010011" when "1000001",
		"00100100110" when "1000010",
		"00110111000" when "1000011",
		"01001001001" when "1000100",
		"01011011000" when "1000101",
		"01101100110" when "1000110",
		"01111110010" when "1000111",
		"10001111100" when "1001000",
		"10100000010" when "1001001",
		"10110000110" when "1001010",
		"11000000110" when "1001011",
		"11010000010" when "1001100",
		"11011111011" when "1001101",
		"11101101111" when "1001110",
		"11111011110" when "1001111",
		"00001001001" when "1010000",
		"00010101110" when "1010001",
		"00100001111" when "1010010",
		"00101101001" when "1010011",
		"00110111110" when "1010100",
		"01000001101" when "1010101",
		"01001010101" when "1010110",
		"01010010111" when "1010111",
		"01011010011" when "1011000",
		"01100001000" when "1011001",
		"01100110110" when "1011010",
		"01101011110" when "1011011",
		"01101111110" when "1011100",
		"01110010111" when "1011101",
		"01110101001" when "1011110",
		"01110110100" when "1011111",
		"01110111000" when "1100000",
		"01110110100" when "1100001",
		"01110101001" when "1100010",
		"01110010111" when "1100011",
		"01101111110" when "1100100",
		"01101011110" when "1100101",
		"01100110110" when "1100110",
		"01100001000" when "1100111",
		"01011010011" when "1101000",
		"01010010111" when "1101001",
		"01001010101" when "1101010",
		"01000001101" when "1101011",
		"00110111110" when "1101100",
		"00101101001" when "1101101",
		"00100001111" when "1101110",
		"00010101110" when "1101111",
		"00001001001" when "1110000",
		"11111011110" when "1110001",
		"11101101111" when "1110010",
		"11011111011" when "1110011",
		"11010000010" when "1110100",
		"11000000110" when "1110101",
		"10110000110" when "1110110",
		"10100000010" when "1110111",
		"10001111100" when "1111000",
		"01111110010" when "1111001",
		"01101100110" when "1111010",
		"01011011000" when "1111011",
		"01001001001" when "1111100",
		"00110111000" when "1111101",
		"00100100110" when "1111110",
		"00010010011" when "1111111",
		"00000000000" when others;
end DataFlow;
