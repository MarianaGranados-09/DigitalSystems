library IEEE;
use IEEE.std_logic_1164.all;

entity ROM_a is 
	port(
		SEL : in std_logic_vector(3 downto 0);
		QOUT : out std_logic_vector(31 downto 0)
		);
end ROM_a;

architecture DataFlow of ROM_a is
begin	
	
	with SEL Select QOUT <=
	"00010000000000000000000000000000" when "0000", --a0
	"11011010110110100011000010101010" when "0001",	--a1
	"00000001001111100111101001111000" when "0010",	--a2
	"00011111110111100001011110001010" when "0011",	--a3
	"00011001100100011011000011111101" when "0100",	--a4
	"11001111010111100110000011001111" when "0101",	--a5
	"11111011000010110110011101101100" when "0110",	--a6
	"00001010110011111101111111111001" when "0111",	--a7	
	"00001101010111010101111100110001" when "1000",	--a8
	"11110111101100111110001111101110" when "1001",	--a9
	"00000000001011001010000110010111" when "1010",	--a10
	"00000000000000000000000000000000" when others;	 
	
end DataFlow;
