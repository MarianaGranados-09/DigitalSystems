library IEEE;
use IEEE.std_logic_1164.all;

entity ROM_b is 
	port(
		SEL : in std_logic_vector(3 downto 0);
		QOUT : out std_logic_vector(31 downto 0)
		);
end ROM_b;

architecture DataFlow of ROM_b is
begin	
	
	with SEL Select QOUT <=
	"00000100100101101000100011100000" when "0000", --b0
	"11111111000110110111001111000110" when "0001",	--b1
	"11101010111000110011100011001100" when "0010",	--b2
	"00000001101000110100001100101100" when "0011",	--b3
	"00101000101100010101001111100100" when "0100",	--b4 
	"00000000000000000000000000000000" when "0101",	--b5
	"11010111010011101010110000011100" when "0110",	--b6
	"11111110010111001011110011010100" when "0111",	--b7
	"00010101000111001100011100110100" when "1000",	--b8
	"00000000111001001000110000111010" when "1001",	--b9
	"11111011011010010111011100100000" when "1010",	--b10
	"00000000000000000000000000000000" when others;	 --b11
	
end DataFlow;
